`timescale 1ns / 1ps

module DECODER(input [31:0] inst,output [4:0] rs2,rd,output reg [4:0] rs1,output reg [63:0] immediate,output reg [3:0] AluFunc,output reg bsel,mwr,werf,type,reg [1:0] wdsel, pcsel);
    wire [6:0] opcode,func7,func6;
    wire [2:0] func3;
    assign rs2 = inst[24:20];
    assign rd = inst[11:7];
    assign opcode = inst[6:0];
    assign func3 = inst[14:12];
    assign func7 = inst[31:25];
    assign func6 = inst[31:26];
//  add, sub, ld, sd, addi, or, and, xor_i,
//  slli, srli, srai
//  jal, jalr    
    
//  bsel -> chooses between the inputs of R-type and I-type to be sent in the ALU
//  wdsel -> take output of MEM or ALU
//  mwr -> MEM write enable
//  werf -> RF write enable
    
    always@(*) begin
        case(opcode)
            7'b0110011 : begin     // R - type
                    if(func3 == 3'b000)begin   
                        if(func7==7'b0000000)
                            AluFunc = 4'b0000;      //ADD   -   add
                        else if(func7==7'b0100000)
                            AluFunc = 4'b0001;      //SUBTRACT -   sub
                    end
                    else if(func3 == 3'b111)begin   //AND   -   and
                        AluFunc = 4'b0010;
                    end
                    else if(func3 == 3'b110)begin   //OR    -   or
                        AluFunc = 4'b0011;
                    end
                    else if(func3 == 3'b100)begin
                        AluFunc = 4'b0100;
                    end
                    bsel=0;
                    wdsel=2'b0;
                    mwr = 0;
                    werf=1;
                    pcsel = 2'b00;
                    type = 1;
                    rs1 = inst[19:15];
            end
            7'b0010011 : begin     //I - type arithmetic
                    if(func3 == 3'b000)begin   
                        AluFunc = 4'b0000;          //ADD_I -   addi
                        immediate = {{52{inst[31]}},inst[31:20]};
                    end
                    else if(func3 == 3'b100)begin   //XOR_I -   xori
                        AluFunc = 4'b0100;
                        immediate = {{52{inst[31]}},inst[31:20]};
                    end
                    else if(func3 == 3'b001)begin
                        if (func6 == 6'b000000)
                            AluFunc = 4'b0101;     //SLL_I -   slli
                        immediate = {{58{inst[31]}},inst[25:20]};
                    end
                    else if(func3 == 3'b101)begin   
                        if(func6 == 6'b000000)
                            AluFunc = 4'b0110;      //SRL_I -   srli
                        else if(func6 == 6'b010000) 
                            AluFunc = 4'b0111;      //SRA_I -   srai
                        immediate = {{58{inst[31]}},inst[25:20]};
                    end
                    bsel = 1;
                    wdsel=0;
                    mwr = 0;
                    werf=1;
                    pcsel = 2'b0;
                    type = 1;
                    rs1 = inst[19:15];
            end
            7'b0000011 : begin     //I - type load
                    if(func3 == 3'b011)begin    //LOAD_DOUBLE   ld
                        AluFunc = 0000;                   
                        type = 1;
                    end
                    if(func3 == 3'b010)begin    //LOAD_WORD   lw
                        AluFunc = 0000;                    
                        type = 0;
                    end
                    bsel = 1;
                    immediate = {{52{inst[31]}},inst[31:20]};
                    wdsel = 1;
                    mwr = 0;
                    werf=1;   
                    pcsel = 2'b0;
                    rs1 = inst[19:15];
            end
            7'b0100011 : begin     //S - type 
                    if(func3 == 3'b111)begin
                        immediate = {{52{inst[31]}},inst[31:26],inst[11:7]};
                        wdsel = 0;
                        bsel=1;
                        AluFunc = 0000;
                        mwr = 1;
                        werf=0;
                        pcsel = 2'b0;                    
                        type = 1;
                        rs1 = inst[19:15];
                    end
            end
            7'b1100011 : begin     //SB - type
                    if(func3 == 3'b000)             // BEQ
                        AluFunc = 4'b1000;
                    else if (func3 == 3'b001)       //BNE
                        AluFunc = 4'b1001;
                    else if (func3 == 3'b100)       //BLT
                        AluFunc = 4'b1010;
                    else if (func3 == 3'b101)       //BGE
                        AluFunc = 4'b1011;
                    immediate = {{52{inst[31]}},inst[7],inst[30:25],inst[11:8],1'b0};
                    wdsel = 0;
                    bsel=0;
                    mwr = 0;
                    werf=0;
                    pcsel = 2'b01;                    
                    type = 1;
                    rs1 = inst[19:15];
            end
            7'b1100111 : begin     //I-type
                    if(func3 == 3'b000)             //JALR
                        AluFunc = 4'b0000;
                    immediate = {{58{inst[31]}},inst[25:20]};
                    wdsel = 2'b10;
                    bsel=1;
                    mwr = 0;
                    werf=1;
                    pcsel = 2'b10;                    
                    type = 1;
                    rs1 = inst[19:15];
            end
            7'b1101111 : begin     //UJ - type
                    AluFunc = 4'b0000;          //JAL
//                    immediate = {{58{inst[31]}},inst[25:20]};
                    immediate = {{44{inst[31]}},inst[19:12],inst[20],inst[30:21],1'b0};
                    wdsel = 2'b10;
                    bsel=1;
                    mwr = 0;
                    werf=1;
                    pcsel = 2'b11;                    
                    type = 1;
                    rs1 = 5'b0;
            end
        endcase
    end
endmodule